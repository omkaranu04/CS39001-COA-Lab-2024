`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/27/2024 05:49:53 PM
// Design Name: 
// Module Name: Instruction_Memory
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module Instruction_Memory #(parameter BRAM_ADDR_WIDTH = 2, BRAM_DATA_WIDTH = 32) (clk, rst, addr, wr_n, rd_n, bram_data_in, bram_data_out);

    input clk, wr_n, rd_n, rst;
    input [BRAM_ADDR_WIDTH-1:0] addr;
    input [BRAM_DATA_WIDTH-1:0] bram_data_in;
    output reg [BRAM_DATA_WIDTH-1:0] bram_data_out;

    reg [BRAM_DATA_WIDTH-1:0] mem [(1<<BRAM_ADDR_WIDTH)-1:0];
    integer i;
//    initial begin
//        // $monitor("ins mem[%d] = %d at %d", 0, mem[0], $time);
//        $readmemb("Instruction_Memory.mem", mem);
//    end

    always @(negedge clk) begin
        // if (wr_n == 1'b0) mem[(addr)] <= bram_data_in;
        if(rst) begin
//            ins for 10 to 1 addition in loop
//            mem[0]=32'b01110100000000010000000000000000; 
//            mem[1]=32'b10010100001000010000000000000100;
//            mem[2]=32'b00000000001000100001000000000000;
//            mem[3]=32'b00001100001000010000000000000001;
//            mem[4]=32'b10011011111111111111111111111101;
//            mem[5]=32'b00011000000000000000000000000000;
            
//            mem[0] = 32'b00000100001000000000000000111100;
//            mem[1] = 32'b01110100000000100000000000000000;
//            mem[2] = 32'b01000100001000010000000000000001;
//            mem[2] = 32'b00011000000000000000000000000000;

// Insertion Sort Instructions

//            mem[0]  = 32'b00000100000000010000000000000001;
//            mem[1]  = 32'b01101100001001000000000000010100;
//            mem[2]  = 32'b10010100100001000000000000001101;
//            mem[3]  = 32'b00001100001000100000000000000001;
//            mem[4]  = 32'b01110100001000110000000000000000;
//            mem[5]  = 32'b10000100010000100000000000000111;
//            mem[6]  = 32'b01110100010001010000000000000000;
//            mem[7]  = 32'b00000000011001010010000000001101;
//            mem[8]  = 32'b10010100100001000000000000000100;
//            mem[9]  = 32'b01111100101000100000000000000001;
//            mem[10] = 32'b00001100010000100000000000000001;
//            mem[11] = 32'b10011011111111111111111111111010;
//            mem[12] = 32'b01111100011000100000000000000001;
//            mem[13] = 32'b00000100001000010000000000000001;
//            mem[14] = 32'b10011011111111111111111111110011;
//            mem[15] = 32'b01110100000000010000000000000000;
//            mem[16] = 32'b01110100000000100000000000000001;
//            mem[17] = 32'b01110100000000110000000000000010;
//            mem[18] = 32'b01110100000001000000000000000011;
//            mem[19] = 32'b01110100000001010000000000000100;
//            mem[20] = 32'b01110100000001100000000000000101;
//            mem[21] = 32'b01110100000001110000000000000110;
//            mem[22] = 32'b01110100000010000000000000000111;
//            mem[23] = 32'b01110100000010010000000000001000;
//            mem[24] = 32'b01110100000010100000000000001001;
//            mem[25] = 32'b00011000000000000000000000000000;

// Booth Algo Working
//            mem[0]  = 32'b00000100000000011111111111110001;
//            mem[1]  = 32'b00000100000000100000000000001110;
//            mem[2]  = 32'b00000100000000110000000000100000;
//            mem[3]  = 32'b00010000011010100101011111111111;
//            mem[4]  = 32'b00001100011010110000000000000001;
//            mem[5]  = 32'b00000100000001000000000000000000;
//            mem[6]  = 32'b00000100000001010000000000000000;
//            mem[7]  = 32'b00010100010001110000000000000001;
//            mem[8]  = 32'b00000000111001010100000000000001;
//            mem[9]  = 32'b10010101000010000000000000000101;
//            mem[10] = 32'b10001101000010000000000000000011;
//            mem[11] = 32'b00000000100000010010011111100000;
//            mem[12] = 32'b10011000000000000000000000000010;
//            mem[13] = 32'b00000000100000010010011111100001;
//            mem[14] = 32'b00010100100001100000000000000001;
//            mem[15] = 32'b01001100100001000000000000000001;
//            mem[16] = 32'b01001100010000100000000000000001;
//            mem[17] = 32'b00000000110010110011000000001000;
//            mem[18] = 32'b00000000010001100001000000000000;
//            mem[19] = 32'b00010000111000000010100000000000;
//            mem[20] = 32'b00001101010010100000000000000001;
//            mem[21] = 32'b10010101010010100000000000000010;
//            mem[22] = 32'b10001101010010101111111111110001;
//            mem[23] = 32'b01000100100001000000000000100000;
//            mem[24] = 32'b00000000010001000001011001100000;
//            mem[25] = 32'b00011000000000000000000000000000;

// CMOV
//            mem[0] = 32'b00000100000000011111111111110100;
//            mem[1] = 32'b00000100000000110000000000000001;
//            mem[2] = 32'b00100000001000110001000000000000;
//            mem[3] = 32'b00000000010000000001000000001111;
//            mem[4] = 32'b00011000000000000000000000000000;

// NON RES DIV
            mem[0]  = 32'b00000100000011100000000000000000;
            mem[1]  = 32'b00000100000000010000000000001111;
            mem[2]  = 32'b01110100000001000000000000000000;
            mem[3]  = 32'b01110100000001010000000000000001;
            mem[4]  = 32'b01000100101001010000000000001111;
            mem[5]  = 32'b01000100100001000000000000000001;
            mem[6]  = 32'b10000100100001000000000000000011;
            mem[7]  = 32'b00000000100001010010000000000001;
            mem[8]  = 32'b10011000000000000000000000000010;
            mem[9]  = 32'b00000000100001010010000000000000;
            mem[10] = 32'b10000100100001000000000000000010;
            mem[11] = 32'b00000100100001000000000000000001;
            mem[12] = 32'b00001100001000010000000000000001;
            mem[13] = 32'b10010100001000010000000000000010;
            mem[14] = 32'b10011011111111111111111111110111;
            mem[15] = 32'b10010100100001000000000000000011;
            mem[16] = 32'b10001100100001000000000000000010;
            mem[17] = 32'b00000000100001010010000000000000;
            mem[18] = 32'b00010100100000100111111111111111;
            mem[19] = 32'b00010100100000111111111111111111;
            mem[20] = 32'b01010100011000110000000000001111;
            mem[21] = 32'b01111100010000000000000000000000;
            mem[22] = 32'b01111100011000000000000000000001;
            mem[23] = 32'b00011000000000000000000000000000;
        end
        else begin
            if (rd_n == 1'b1) bram_data_out <= mem[addr];
        end 
    end

endmodule

